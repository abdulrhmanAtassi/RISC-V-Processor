module hazard_unit (
    input [4:0] id_ex_rs, id_ex_rt, ex_mem_rd, mem_wb_rd,
    input ex_mem_reg_write, mem_wb_reg_write,
    output stall
);
    // Hazard detection logic goes here
endmodule
