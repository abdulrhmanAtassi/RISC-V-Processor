module if_stage (
    input clk,
    input reset,
    input [31:0] pc_in,
    output [31:0] pc_out,
    output [31:0] instruction
);
    // IF stage logic goes here
endmodule
